assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i) |-> i2c_master_top.wb_ack_o);:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && !i2c_master_top.wb_ack_o) |-> ##1 i2c_master_top.wb_ack_o);
assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_we_i |-> i2c_master_top.wb_wacc);:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_we_i && i2c_master_top.wb_ack_o) |-> i2c_master_top.wb_wacc);
assert property (@(posedge i2c_master_top.wb_clk_i)!i2c_master_top.wb_stb_i |-> !i2c_master_top.wb_ack_o);:assert property (@(posedge i2c_master_top.wb_clk_i)!i2c_master_top.wb_stb_i |-> ##1 !i2c_master_top.wb_ack_o);
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b000 |-> ##1 i2c_master_top.wb_dat_o == i2c_master_top.prer[7:0]);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b000 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[7:0]));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b010 |-> ##1 i2c_master_top.wb_dat_o == i2c_master_top.ctr);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b010 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.ctr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b010 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b011 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b101 |-> i2c_master_top.wb_dat_o == $past(i2c_master_top.sr));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b100 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.sr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b101 |-> i2c_master_top.wb_dat_o == $past(i2c_master_top.txr));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b101 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.txr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b110 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b011 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b111 |-> ##1 i2c_master_top.wb_dat_o == 1);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b111 |-> ##1 i2c_master_top.wb_dat_o == 0);
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i |-> (i2c_master_top.wb_dat_o[0] == 0 || i2c_master_top.wb_dat_o[0] == 0));:assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i |-> (i2c_master_top.wb_dat_o[0] == 1 || i2c_master_top.wb_dat_o[0] == 0));
assert property (@(posedge i2c_master_top.wb_clk_i)(i2c_master_top.wb_adr_i == 3'b000 || i2c_master_top.wb_adr_i == 3'b001 || i2c_master_top.wb_adr_i == 3'b010 ||i2c_master_top.wb_adr_i == 3'b011 || i2c_master_top.wb_adr_i == 3'b100 || i2c_master_top.wb_adr_i == 3'b101 ||i2c_master_top.wb_adr_i == 3'b110 || i2c_master_top.wb_adr_i == 3'b111)|-> ##1 (i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[7:0]) || i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[15:8]) || i2c_master_top.wb_dat_o == i2c_master_top.ctr || i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr) || i2c_master_top.wb_dat_o == $past(i2c_master_top.sr) || i2c_master_top.wb_dat_o == i2c_master_top.txr || i2c_master_top.wb_dat_o == $past(i2c_master_top.cr) || i2c_master_top.wb_dat_o == 0));:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_adr_i == 3'b000 || i2c_master_top.wb_adr_i == 3'b001 || i2c_master_top.wb_adr_i == 3'b010 || i2c_master_top.wb_adr_i == 3'b011 || i2c_master_top.wb_adr_i == 3'b100 || i2c_master_top.wb_adr_i == 3'b101 || i2c_master_top.wb_adr_i == 3'b110 || i2c_master_top.wb_adr_i == 3'b111)|-> ##1 (i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[7:0]) || i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[15:8]) || i2c_master_top.wb_dat_o == $past(i2c_master_top.ctr) || i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr) || i2c_master_top.wb_dat_o == $past(i2c_master_top.sr) || i2c_master_top.wb_dat_o == $past(i2c_master_top.txr) || i2c_master_top.wb_dat_o == $past(i2c_master_top.cr) || i2c_master_top.wb_dat_o == 0));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b111 |-> ##1 i2c_master_top.wb_dat_o == 1);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b111 |-> ##1 i2c_master_top.wb_dat_o == 0);
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b000 |-> ##1 i2c_master_top.wb_dat_o == i2c_master_top.prer[7:0]);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b000 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[7:0]));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b001 |-> i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[15:8]));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b001 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.prer[15:8]));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b011 |-> ##2 i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b011 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.rxr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b100 |-> i2c_master_top.wb_dat_o == $past(i2c_master_top.sr));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b100 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.sr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b100 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.txr));:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b101 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.txr));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_adr_i == 3'b110 |-> ##1 i2c_master_top.wb_dat_o == i2c_master_top.cr);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_adr_i == 3'b110 |-> ##1 i2c_master_top.wb_dat_o == $past(i2c_master_top.cr));
assert property (@(posedge i2c_master_top.wb_clk_i)(i2c_master_top.wb_adr_i == 3'b000) |-> (i2c_master_top.wb_adr_i == 3'b001 || i2c_master_top.wb_adr_i == 3'b010 || i2c_master_top.wb_adr_i == 3'b100 || i2c_master_top.wb_adr_i == 3'b101 || i2c_master_top.wb_adr_i == 3'b110));:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_adr_i == 3'b000) |-> !(i2c_master_top.wb_adr_i == 3'b001 || i2c_master_top.wb_adr_i == 3'b010 || i2c_master_top.wb_adr_i == 3'b011 || i2c_master_top.wb_adr_i == 3'b100 || i2c_master_top.wb_adr_i == 3'b101 || i2c_master_top.wb_adr_i == 3'b110));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.core_en && i2c_master_top.wb_adr_i == 3'b101 |-> i2c_master_top.cr == i2c_master_top.wb_dat_i);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.core_en && i2c_master_top.wb_adr_i == 3'b100 |-> i2c_master_top.cr == i2c_master_top.wb_dat_i);
assert property (@(posedge i2c_master_bit_ctrl.clk) disable iff(i2c_master_bit_ctrl.nReset) i2c_master_bit_ctrl.nReset || i2c_master_bit_ctrl.rst |-> ##1 i2c_master_bit_ctrl.cSCL == 2'b00);:assert property (@(posedge i2c_master_bit_ctrl.clk) !i2c_master_bit_ctrl.nReset || i2c_master_bit_ctrl.rst |-> ##1 i2c_master_bit_ctrl.cSCL == 2'b00);
assert property (@(posedge i2c_master_bit_ctrl.clk)!i2c_master_bit_ctrl.nReset || !i2c_master_bit_ctrl.rst |-> i2c_master_bit_ctrl.cSDA == 2'b00);:assert property (@(posedge i2c_master_bit_ctrl.clk) !i2c_master_bit_ctrl.nReset || i2c_master_bit_ctrl.rst |-> ##1 i2c_master_bit_ctrl.cSDA == 2'b00);
assert property (@(posedge i2c_master_top.wb_clk_i) (!i2c_master_top.rst_i == (i2c_master_top.arst_i ^ i2c_master_top.ARST_LVL)));:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.rst_i == (i2c_master_top.arst_i ^ i2c_master_top.ARST_LVL)));
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_wacc |-> !i2c_master_top.wb_we_i);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_wacc |-> i2c_master_top.wb_we_i);//下面的波形图可能要重新收集
assert property (@(posedge i2c_master_top.wb_clk_i)i2c_master_top.wb_cyc_i |-> ##1 (i2c_master_top.wb_ack_o == 1'b0));:assert property (@(posedge i2c_master_top.wb_clk_i) (!i2c_master_top.wb_cyc_i || !i2c_master_top.wb_stb_i) |-> ##1 (i2c_master_top.wb_ack_o == 1'b0));
assert property (@(posedge i2c_master_top.wb_clk_i)($past(i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i) && (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i)) |-> (i2c_master_top.wb_ack_o != $past(i2c_master_top.wb_ack_o)));:assert property (@(posedge i2c_master_top.wb_clk_i) ($past(i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i) && (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i)) |=> (i2c_master_top.wb_ack_o != $past(i2c_master_top.wb_ack_o)));
assert property (@(posedge i2c_master_top.wb_clk_i)(i2c_master_top.ien == 1'b0) |-> (i2c_master_top.wb_inta_o == 1'b0));:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.ien == 1'b0) |=> (i2c_master_top.wb_inta_o == 1'b0));
assert property (@(posedge i2c_master_top.wb_clk_i) disable iff (!i2c_master_top.rst_i)i2c_master_top.ctr[7] == 1'b0 |-> i2c_master_top.byte_controller.ena == 1'b1);:assert property (@(posedge i2c_master_top.wb_clk_i) disable iff (!i2c_master_top.rst_i) i2c_master_top.ctr[7] == 1'b1 |-> i2c_master_top.byte_controller.ena == 1'b1);
assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_rst_i == 1'b1) |->(i2c_master_top.ctr == 8'h00));:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.rst_i == 1'b0) |->(i2c_master_top.ctr == 8'h00));
assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_rst_i |-> !i2c_master_top.cr);:assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.rst_i==1'b0 |-> !i2c_master_top.cr);
assert property (@(posedge i2c_master_top.wb_clk_i) i2c_master_top.wb_rst_i |-> !i2c_master_top.tip);:assert property (@(posedge i2c_master_top.wb_clk_i) !i2c_master_top.rst_i |-> !i2c_master_top.tip);
assert property  (@(posedge i2c_master_top.wb_clk_i) disable iff (!i2c_master_top.wb_rst_i) (i2c_master_top.wb_stb_i && i2c_master_top.wb_cyc_i) |-> ((i2c_master_top.wb_adr_i >= 3'b000) && (i2c_master_top.wb_adr_i <= 3'b100)));:assert property  (@(posedge i2c_master_top.wb_clk_i) disable iff (!i2c_master_top.wb_rst_i) (i2c_master_top.wb_adr_i >= 3'b000) && (i2c_master_top.wb_adr_i <= 3'b100));
assert property  (@(posedge i2c_master_top.wb_clk_i) disable iff (!i2c_master_top.wb_rst_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && !i2c_master_top.wb_we_i) |-> !($isunknown(i2c_master_top.wb_dat_o)));:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && !i2c_master_top.wb_ack_o) |-> ##1 i2c_master_top.wb_ack_o);
assert property  (@(posedge i2c_master_top.wb_clk_i) disable iff (i2c_master_top.wb_rst_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && i2c_master_top.wb_we_i) |-> i2c_master_top.wb_adr_i == 0);:assert property  (@(posedge i2c_master_top.wb_clk_i) disable iff (i2c_master_top.wb_rst_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && i2c_master_top.wb_we_i) |-> $isunknown(i2c_master_top.wb_adr_i) == 0 && $isunknown(i2c_master_top.wb_dat_i) == 0);
assert property  (@(posedge i2c_master_top.wb_clk_i) disable iff (i2c_master_top.wb_rst_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && i2c_master_top.wb_we_i) |=> ##[1:2] i2c_master_top.wb_ack_o);:assert property (@(posedge i2c_master_top.wb_clk_i) (i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && !i2c_master_top.wb_ack_o) |-> ##[1:2] i2c_master_top.wb_ack_o);
assert property  (@(posedge i2c_master_top.wb_clk_i) !i2c_master_top.rst_i |-> !(i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && i2c_master_top.wb_we_i));:assert property  (@(posedge i2c_master_top.wb_clk_i) !i2c_master_top.rst_i |-> ##1 !(i2c_master_top.wb_cyc_i && i2c_master_top.wb_stb_i && i2c_master_top.wb_we_i));













